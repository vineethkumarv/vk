package pack1;
  function test;
    $display("hi this this is pack1");
  endfunction
endpackage
