module one;
int a;
string k;
initial begin
    if(type(type(k))==type(int)) $display(/*"%0s",type(k)*/"string");
    $display(k);
  end
  endmodule

